----------------------------------------------------------------------------------
-- Engineer: Diego Ceresuela, Oscar Clemente.
-- 
-- Create Date: 13.04.2016 08:23:25
-- Module Name: sigmoid - Behavioral
-- Description: Implements a ROM containing the aproximation of the sigmoid function.
-- 
-- Dependencies: 
-- 
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sigmoid is
    Port ( Y : in STD_LOGIC_VECTOR (31 downto 0);
           O : out STD_LOGIC_VECTOR (31 downto 0);
           clk: in STD_LOGIC );
end sigmoid;

architecture Behavioral of sigmoid is

type rom is array (0 to 3410) of STD_LOGIC_VECTOR (15 downto 0);
    signal sigmoid_val : rom := (x"0000",x"0001",x"0001",x"0001",x"0001",x"0001",x"0002",x"0002",x"0003",x"0003",x"0003",x"0003",x"0003",x"0003",x"0004",x"0004",x"0004",x"0004",x"0004",x"0004",x"0005",x"0005",x"0005",x"0005",x"0006",x"0006",x"0006",x"0007",x"0007",x"0007",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0008",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"0009",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000a",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000b",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000c",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000d",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000e",x"000f",x"000f",x"000f",x"000f",x"000f",x"000f",x"000f",x"000f",x"000f",x"000f",x"000f",x"000f",x"0010",x"0010",x"0010",x"0010",x"0010",x"0010",x"0010",x"0010",x"0010",x"0010",x"0010",x"0011",x"0011",x"0011",x"0011",x"0011",x"0011",x"0011",x"0011",x"0011",x"0011",x"0012",x"0012",x"0012",x"0012",x"0012",x"0012",x"0012",x"0012",x"0012",x"0012",x"0012",x"0013",x"0013",x"0013",x"0013",x"0013",x"0013",x"0013",x"0013",x"0013",x"0014",x"0014",x"0014",x"0014",x"0014",x"0014",x"0014",x"0014",x"0014",x"0015",x"0015",x"0015",x"0015",x"0015",x"0015",x"0015",x"0015",x"0015",x"0016",x"0016",x"0016",x"0016",x"0016",x"0016",x"0016",x"0016",x"0017",x"0017",x"0017",x"0017",x"0017",x"0017",x"0017",x"0017",x"0018",x"0018",x"0018",x"0018",x"0018",x"0018",x"0018",x"0018",x"0019",x"0019",x"0019",x"0019",x"0019",x"0019",x"0019",x"001a",x"001a",x"001a",x"001a",x"001a",x"001a",x"001a",x"001b",x"001b",x"001b",x"001b",x"001b",x"001b",x"001b",x"001c",x"001c",x"001c",x"001c",x"001c",x"001c",x"001d",x"001d",x"001d",x"001d",x"001d",x"001d",x"001d",x"001e",x"001e",x"001e",x"001e",x"001e",x"001e",x"001f",x"001f",x"001f",x"001f",x"001f",x"001f",x"0020",x"0020",x"0020",x"0020",x"0020",x"0021",x"0021",x"0021",x"0021",x"0021",x"0021",x"0022",x"0022",x"0022",x"0022",x"0022",x"0023",x"0023",x"0023",x"0023",x"0023",x"0023",x"0024",x"0024",x"0024",x"0024",x"0024",x"0025",x"0025",x"0025",x"0025",x"0025",x"0026",x"0026",x"0026",x"0026",x"0026",x"0027",x"0027",x"0027",x"0027",x"0028",x"0028",x"0028",x"0028",x"0028",x"0029",x"0029",x"0029",x"0029",x"002a",x"002a",x"002a",x"002a",x"002a",x"002b",x"002b",x"002b",x"002b",x"002c",x"002c",x"002c",x"002c",x"002d",x"002d",x"002d",x"002d",x"002e",x"002e",x"002e",x"002e",x"002f",x"002f",x"002f",x"002f",x"0030",x"0030",x"0030",x"0030",x"0031",x"0031",x"0031",x"0031",x"0032",x"0032",x"0032",x"0033",x"0033",x"0033",x"0033",x"0034",x"0034",x"0034",x"0034",x"0035",x"0035",x"0035",x"0036",x"0036",x"0036",x"0036",x"0037",x"0037",x"0037",x"0038",x"0038",x"0038",x"0039",x"0039",x"0039",x"003a",x"003a",x"003a",x"003a",x"003b",x"003b",x"003b",x"003c",x"003c",x"003c",x"003d",x"003d",x"003d",x"003e",x"003e",x"003e",x"003f",x"003f",x"003f",x"0040",x"0040",x"0040",x"0041",x"0041",x"0041",x"0042",x"0042",x"0043",x"0043",x"0043",x"0044",x"0044",x"0044",x"0045",x"0045",x"0045",x"0046",x"0046",x"0047",x"0047",x"0047",x"0048",x"0048",x"0049",x"0049",x"0049",x"004a",x"004a",x"004b",x"004b",x"004b",x"004c",x"004c",x"004d",x"004d",x"004d",x"004e",x"004e",x"004f",x"004f",x"0050",x"0050",x"0050",x"0051",x"0051",x"0052",x"0052",x"0053",x"0053",x"0054",x"0054",x"0054",x"0055",x"0055",x"0056",x"0056",x"0057",x"0057",x"0058",x"0058",x"0059",x"0059",x"005a",x"005a",x"005b",x"005b",x"005c",x"005c",x"005d",x"005d",x"005e",x"005e",x"005f",x"005f",x"0060",x"0060",x"0061",x"0061",x"0062",x"0062",x"0063",x"0063",x"0064",x"0064",x"0065",x"0065",x"0066",x"0066",x"0067",x"0068",x"0068",x"0069",x"0069",x"006a",x"006a",x"006b",x"006c",x"006c",x"006d",x"006d",x"006e",x"006f",x"006f",x"0070",x"0070",x"0071",x"0072",x"0072",x"0073",x"0073",x"0074",x"0075",x"0075",x"0076",x"0077",x"0077",x"0078",x"0078",x"0079",x"007a",x"007a",x"007b",x"007c",x"007c",x"007d",x"007e",x"007e",x"007f",x"0080",x"0081",x"0081",x"0082",x"0083",x"0083",x"0084",x"0085",x"0085",x"0086",x"0087",x"0088",x"0088",x"0089",x"008a",x"008b",x"008b",x"008c",x"008d",x"008e",x"008e",x"008f",x"0090",x"0091",x"0091",x"0092",x"0093",x"0094",x"0095",x"0095",x"0096",x"0097",x"0098",x"0099",x"0099",x"009a",x"009b",x"009c",x"009d",x"009e",x"009e",x"009f",x"00a0",x"00a1",x"00a2",x"00a3",x"00a4",x"00a5",x"00a5",x"00a6",x"00a7",x"00a8",x"00a9",x"00aa",x"00ab",x"00ac",x"00ad",x"00ae",x"00af",x"00b0",x"00b0",x"00b1",x"00b2",x"00b3",x"00b4",x"00b5",x"00b6",x"00b7",x"00b8",x"00b9",x"00ba",x"00bb",x"00bc",x"00bd",x"00be",x"00bf",x"00c0",x"00c1",x"00c2",x"00c3",x"00c4",x"00c6",x"00c7",x"00c8",x"00c9",x"00ca",x"00cb",x"00cc",x"00cd",x"00ce",x"00cf",x"00d0",x"00d2",x"00d3",x"00d4",x"00d5",x"00d6",x"00d7",x"00d8",x"00da",x"00db",x"00dc",x"00dd",x"00de",x"00df",x"00e1",x"00e2",x"00e3",x"00e4",x"00e6",x"00e7",x"00e8",x"00e9",x"00eb",x"00ec",x"00ed",x"00ee",x"00f0",x"00f1",x"00f2",x"00f4",x"00f5",x"00f6",x"00f7",x"00f9",x"00fa",x"00fb",x"00fd",x"00fe",x"0100",x"0101",x"0102",x"0104",x"0105",x"0107",x"0108",x"0109",x"010b",x"010c",x"010e",x"010f",x"0111",x"0112",x"0113",x"0115",x"0116",x"0118",x"0119",x"011b",x"011c",x"011e",x"0120",x"0121",x"0123",x"0124",x"0126",x"0127",x"0129",x"012b",x"012c",x"012e",x"012f",x"0131",x"0133",x"0134",x"0136",x"0138",x"0139",x"013b",x"013d",x"013e",x"0140",x"0142",x"0143",x"0145",x"0147",x"0149",x"014a",x"014c",x"014e",x"0150",x"0152",x"0153",x"0155",x"0157",x"0159",x"015b",x"015d",x"015f",x"0160",x"0162",x"0164",x"0166",x"0168",x"016a",x"016c",x"016e",x"0170",x"0172",x"0174",x"0176",x"0178",x"017a",x"017c",x"017e",x"0180",x"0182",x"0184",x"0186",x"0188",x"018a",x"018c",x"018f",x"0191",x"0193",x"0195",x"0197",x"0199",x"019c",x"019e",x"01a0",x"01a2",x"01a4",x"01a7",x"01a9",x"01ab",x"01ad",x"01b0",x"01b2",x"01b4",x"01b7",x"01b9",x"01bb",x"01be",x"01c0",x"01c3",x"01c5",x"01c7",x"01ca",x"01cc",x"01cf",x"01d1",x"01d4",x"01d6",x"01d9",x"01db",x"01de",x"01e0",x"01e3",x"01e6",x"01e8",x"01eb",x"01ed",x"01f0",x"01f3",x"01f5",x"01f8",x"01fb",x"01fd",x"0200",x"0203",x"0206",x"0208",x"020b",x"020e",x"0211",x"0214",x"0217",x"0219",x"021c",x"021f",x"0222",x"0225",x"0228",x"022b",x"022e",x"0231",x"0234",x"0237",x"023a",x"023d",x"0240",x"0243",x"0246",x"0249",x"024c",x"0250",x"0253",x"0256",x"0259",x"025c",x"025f",x"0263",x"0266",x"0269",x"026d",x"0270",x"0273",x"0277",x"027a",x"027d",x"0281",x"0284",x"0288",x"028b",x"028e",x"0292",x"0295",x"0299",x"029d",x"02a0",x"02a4",x"02a7",x"02ab",x"02af",x"02b2",x"02b6",x"02ba",x"02bd",x"02c1",x"02c5",x"02c9",x"02cc",x"02d0",x"02d4",x"02d8",x"02dc",x"02e0",x"02e4",x"02e8",x"02ec",x"02f0",x"02f4",x"02f8",x"02fc",x"0300",x"0304",x"0308",x"030c",x"0310",x"0314",x"0319",x"031d",x"0321",x"0325",x"032a",x"032e",x"0332",x"0337",x"033b",x"033f",x"0344",x"0348",x"034d",x"0351",x"0356",x"035a",x"035f",x"0363",x"0368",x"036d",x"0371",x"0376",x"037b",x"037f",x"0384",x"0389",x"038e",x"0393",x"0397",x"039c",x"03a1",x"03a6",x"03ab",x"03b0",x"03b5",x"03ba",x"03bf",x"03c4",x"03c9",x"03cf",x"03d4",x"03d9",x"03de",x"03e3",x"03e9",x"03ee",x"03f3",x"03f9",x"03fe",x"0404",x"0409",x"040e",x"0414",x"0419",x"041f",x"0425",x"042a",x"0430",x"0436",x"043b",x"0441",x"0447",x"044d",x"0452",x"0458",x"045e",x"0464",x"046a",x"0470",x"0476",x"047c",x"0482",x"0488",x"048e",x"0495",x"049b",x"04a1",x"04a7",x"04ae",x"04b4",x"04ba",x"04c1",x"04c7",x"04ce",x"04d4",x"04db",x"04e1",x"04e8",x"04ee",x"04f5",x"04fc",x"0503",x"0509",x"0510",x"0517",x"051e",x"0525",x"052c",x"0533",x"053a",x"0541",x"0548",x"054f",x"0556",x"055d",x"0565",x"056c",x"0573",x"057b",x"0582",x"0589",x"0591",x"0598",x"05a0",x"05a8",x"05af",x"05b7",x"05bf",x"05c6",x"05ce",x"05d6",x"05de",x"05e6",x"05ee",x"05f6",x"05fe",x"0606",x"060e",x"0616",x"061e",x"0626",x"062f",x"0637",x"063f",x"0648",x"0650",x"0659",x"0661",x"066a",x"0672",x"067b",x"0684",x"068d",x"0695",x"069e",x"06a7",x"06b0",x"06b9",x"06c2",x"06cb",x"06d4",x"06dd",x"06e7",x"06f0",x"06f9",x"0702",x"070c",x"0715",x"071f",x"0728",x"0732",x"073c",x"0745",x"074f",x"0759",x"0763",x"076d",x"0777",x"0781",x"078b",x"0795",x"079f",x"07a9",x"07b3",x"07be",x"07c8",x"07d2",x"07dd",x"07e7",x"07f2",x"07fc",x"0807",x"0812",x"081d",x"0827",x"0832",x"083d",x"0848",x"0853",x"085e",x"086a",x"0875",x"0880",x"088b",x"0897",x"08a2",x"08ae",x"08b9",x"08c5",x"08d1",x"08dc",x"08e8",x"08f4",x"0900",x"090c",x"0918",x"0924",x"0930",x"093c",x"0949",x"0955",x"0961",x"096e",x"097a",x"0987",x"0994",x"09a0",x"09ad",x"09ba",x"09c7",x"09d4",x"09e1",x"09ee",x"09fb",x"0a08",x"0a15",x"0a23",x"0a30",x"0a3e",x"0a4b",x"0a59",x"0a67",x"0a74",x"0a82",x"0a90",x"0a9e",x"0aac",x"0aba",x"0ac8",x"0ad7",x"0ae5",x"0af3",x"0b02",x"0b10",x"0b1f",x"0b2d",x"0b3c",x"0b4b",x"0b5a",x"0b69",x"0b78",x"0b87",x"0b96",x"0ba5",x"0bb5",x"0bc4",x"0bd4",x"0be3",x"0bf3",x"0c03",x"0c12",x"0c22",x"0c32",x"0c42",x"0c52",x"0c62",x"0c73",x"0c83",x"0c93",x"0ca4",x"0cb4",x"0cc5",x"0cd6",x"0ce7",x"0cf7",x"0d08",x"0d19",x"0d2b",x"0d3c",x"0d4d",x"0d5e",x"0d70",x"0d82",x"0d93",x"0da5",x"0db7",x"0dc9",x"0ddb",x"0ded",x"0dff",x"0e11",x"0e23",x"0e36",x"0e48",x"0e5b",x"0e6d",x"0e80",x"0e93",x"0ea6",x"0eb9",x"0ecc",x"0edf",x"0ef3",x"0f06",x"0f1a",x"0f2d",x"0f41",x"0f55",x"0f69",x"0f7d",x"0f91",x"0fa5",x"0fb9",x"0fcd",x"0fe2",x"0ff6",x"100b",x"1020",x"1034",x"1049",x"105e",x"1074",x"1089",x"109e",x"10b3",x"10c9",x"10df",x"10f4",x"110a",x"1120",x"1136",x"114c",x"1162",x"1179",x"118f",x"11a6",x"11bc",x"11d3",x"11ea",x"1201",x"1218",x"122f",x"1247",x"125e",x"1275",x"128d",x"12a5",x"12bd",x"12d5",x"12ed",x"1305",x"131d",x"1335",x"134e",x"1366",x"137f",x"1398",x"13b1",x"13ca",x"13e3",x"13fc",x"1416",x"142f",x"1449",x"1463",x"147d",x"1497",x"14b1",x"14cb",x"14e5",x"1500",x"151a",x"1535",x"1550",x"156b",x"1586",x"15a1",x"15bc",x"15d7",x"15f3",x"160f",x"162a",x"1646",x"1662",x"167f",x"169b",x"16b7",x"16d4",x"16f0",x"170d",x"172a",x"1747",x"1764",x"1782",x"179f",x"17bd",x"17da",x"17f8",x"1816",x"1834",x"1852",x"1871",x"188f",x"18ae",x"18cc",x"18eb",x"190a",x"1929",x"1949",x"1968",x"1988",x"19a7",x"19c7",x"19e7",x"1a07",x"1a27",x"1a48",x"1a68",x"1a89",x"1aaa",x"1aca",x"1aec",x"1b0d",x"1b2e",x"1b50",x"1b71",x"1b93",x"1bb5",x"1bd7",x"1bf9",x"1c1b",x"1c3e",x"1c61",x"1c83",x"1ca6",x"1cc9",x"1cec",x"1d10",x"1d33",x"1d57",x"1d7b",x"1d9f",x"1dc3",x"1de7",x"1e0b",x"1e30",x"1e55",x"1e79",x"1e9e",x"1ec4",x"1ee9",x"1f0e",x"1f34",x"1f5a",x"1f80",x"1fa6",x"1fcc",x"1ff2",x"2019",x"203f",x"2066",x"208d",x"20b4",x"20dc",x"2103",x"212b",x"2153",x"217b",x"21a3",x"21cb",x"21f3",x"221c",x"2245",x"226e",x"2297",x"22c0",x"22e9",x"2313",x"233c",x"2366",x"2390",x"23ba",x"23e5",x"240f",x"243a",x"2465",x"2490",x"24bb",x"24e6",x"2512",x"253e",x"2569",x"2595",x"25c2",x"25ee",x"261a",x"2647",x"2674",x"26a1",x"26ce",x"26fc",x"2729",x"2757",x"2785",x"27b3",x"27e1",x"280f",x"283e",x"286d",x"289b",x"28cb",x"28fa",x"2929",x"2959",x"2988",x"29b8",x"29e9",x"2a19",x"2a49",x"2a7a",x"2aab",x"2adc",x"2b0d",x"2b3e",x"2b70",x"2ba1",x"2bd3",x"2c05",x"2c37",x"2c6a",x"2c9c",x"2ccf",x"2d02",x"2d35",x"2d68",x"2d9c",x"2dd0",x"2e03",x"2e37",x"2e6b",x"2ea0",x"2ed4",x"2f09",x"2f3e",x"2f73",x"2fa8",x"2fde",x"3013",x"3049",x"307f",x"30b5",x"30eb",x"3122",x"3159",x"3190",x"31c7",x"31fe",x"3235",x"326d",x"32a5",x"32dc",x"3315",x"334d",x"3385",x"33be",x"33f7",x"3430",x"3469",x"34a3",x"34dc",x"3516",x"3550",x"358a",x"35c4",x"35ff",x"363a",x"3674",x"36af",x"36eb",x"3726",x"3762",x"379d",x"37d9",x"3816",x"3852",x"388e",x"38cb",x"3908",x"3945",x"3982",x"39c0",x"39fd",x"3a3b",x"3a79",x"3ab7",x"3af5",x"3b34",x"3b72",x"3bb1",x"3bf0",x"3c30",x"3c6f",x"3cae",x"3cee",x"3d2e",x"3d6e",x"3daf",x"3def",x"3e30",x"3e70",x"3eb1",x"3ef3",x"3f34",x"3f76",x"3fb7",x"3ff9",x"403b",x"407e",x"40c0",x"4103",x"4145",x"4188",x"41cb",x"420f",x"4252",x"4296",x"42da",x"431e",x"4362",x"43a6",x"43eb",x"442f",x"4474",x"44b9",x"44ff",x"4544",x"458a",x"45cf",x"4615",x"465b",x"46a1",x"46e8",x"472e",x"4775",x"47bc",x"4803",x"484a",x"4892",x"48d9",x"4921",x"4969",x"49b1",x"49f9",x"4a42",x"4a8a",x"4ad3",x"4b1c",x"4b65",x"4bae",x"4bf8",x"4c41",x"4c8b",x"4cd5",x"4d1f",x"4d69",x"4db3",x"4dfe",x"4e48",x"4e93",x"4ede",x"4f29",x"4f75",x"4fc0",x"500c",x"5057",x"50a3",x"50ef",x"513b",x"5188",x"51d4",x"5221",x"526e",x"52ba",x"5308",x"5355",x"53a2",x"53f0",x"543d",x"548b",x"54d9",x"5527",x"5575",x"55c4",x"5612",x"5661",x"56af",x"56fe",x"574d",x"579d",x"57ec",x"583b",x"588b",x"58db",x"592a",x"597a",x"59ca",x"5a1b",x"5a6b",x"5abc",x"5b0c",x"5b5d",x"5bae",x"5bff",x"5c50",x"5ca1",x"5cf2",x"5d44",x"5d95",x"5de7",x"5e39",x"5e8b",x"5edd",x"5f2f",x"5f81",x"5fd4",x"6026",x"6079",x"60cc",x"611e",x"6171",x"61c4",x"6217",x"626b",x"62be",x"6312",x"6365",x"63b9",x"640c",x"6460",x"64b4",x"6508",x"655c",x"65b1",x"6605",x"6659",x"66ae",x"6703",x"6757",x"67ac",x"6801",x"6856",x"68ab",x"6900",x"6955",x"69ab",x"6a00",x"6a55",x"6aab",x"6b00",x"6b56",x"6bac",x"6c02",x"6c58",x"6cad",x"6d04",x"6d5a",x"6db0",x"6e06",x"6e5c",x"6eb3",x"6f09",x"6f60",x"6fb6",x"700d",x"7063",x"70ba",x"7111",x"7168",x"71bf",x"7216",x"726d",x"72c4",x"731b",x"7372",x"73c9",x"7420",x"7477",x"74cf",x"7526",x"757d",x"75d5",x"762c",x"7684",x"76db",x"7733",x"778b",x"77e2",x"783a",x"7892",x"78e9",x"7941",x"7999",x"79f1",x"7a48",x"7aa0",x"7af8",x"7b50",x"7ba8",x"7c00",x"7c58",x"7cb0",x"7d08",x"7d60",x"7db7",x"7e0f",x"7e67",x"7ebf",x"7f17",x"7f6f",x"7fc7",x"801f",x"8077",x"80cf",x"8127",x"817f",x"81d7",x"822f",x"8287",x"82df",x"8337",x"838f",x"83e7",x"843f",x"8497",x"84ef",x"8547",x"859e",x"85f6",x"864e",x"86a6",x"86fe",x"8755",x"87ad",x"8805",x"885c",x"88b4",x"890c",x"8963",x"89bb",x"8a12",x"8a6a",x"8ac1",x"8b18",x"8b70",x"8bc7",x"8c1e",x"8c75",x"8ccc",x"8d24",x"8d7b",x"8dd2",x"8e29",x"8e7f",x"8ed6",x"8f2d",x"8f84",x"8fda",x"9031",x"9088",x"90de",x"9135",x"918b",x"91e1",x"9238",x"928e",x"92e4",x"933a",x"9390",x"93e6",x"943c",x"9491",x"94e7",x"953d",x"9592",x"95e8",x"963d",x"9692",x"96e8",x"973d",x"9792",x"97e7",x"983c",x"9890",x"98e5",x"993a",x"998e",x"99e3",x"9a37",x"9a8b",x"9ae0",x"9b34",x"9b88",x"9bdb",x"9c2f",x"9c83",x"9cd7",x"9d2a",x"9d7d",x"9dd1",x"9e24",x"9e77",x"9eca",x"9f1d",x"9f6f",x"9fc2",x"a015",x"a067",x"a0b9",x"a10c",x"a15e",x"a1b0",x"a201",x"a253",x"a2a5",x"a2f6",x"a348",x"a399",x"a3ea",x"a43b",x"a48c",x"a4dd",x"a52d",x"a57e",x"a5ce",x"a61e",x"a66f",x"a6bf",x"a70e",x"a75e",x"a7ae",x"a7fd",x"a84d",x"a89c",x"a8eb",x"a93a",x"a989",x"a9d7",x"aa26",x"aa74",x"aac2",x"ab11",x"ab5f",x"abac",x"abfa",x"ac48",x"ac95",x"ace2",x"ad2f",x"ad7c",x"adc9",x"ae16",x"ae62",x"aeaf",x"aefb",x"af47",x"af93",x"afdf",x"b02a",x"b076",x"b0c1",x"b10c",x"b157",x"b1a2",x"b1ed",x"b237",x"b282",x"b2cc",x"b316",x"b360",x"b3aa",x"b3f3",x"b43d",x"b486",x"b4cf",x"b518",x"b561",x"b5a9",x"b5f2",x"b63a",x"b682",x"b6ca",x"b712",x"b75a",x"b7a1",x"b7e8",x"b82f",x"b876",x"b8bd",x"b904",x"b94a",x"b991",x"b9d7",x"ba1d",x"ba62",x"baa8",x"baed",x"bb33",x"bb78",x"bbbd",x"bc01",x"bc46",x"bc8a",x"bccf",x"bd13",x"bd57",x"bd9a",x"bdde",x"be21",x"be64",x"bea7",x"beea",x"bf2d",x"bf6f",x"bfb2",x"bff4",x"c036",x"c077",x"c0b9",x"c0fa",x"c13c",x"c17d",x"c1be",x"c1fe",x"c23f",x"c27f",x"c2bf",x"c2ff",x"c33f",x"c37f",x"c3be",x"c3fd",x"c43c",x"c47b",x"c4ba",x"c4f9",x"c537",x"c575",x"c5b3",x"c5f1",x"c62f",x"c66c",x"c6a9",x"c6e6",x"c723",x"c760",x"c79d",x"c7d9",x"c815",x"c851",x"c88d",x"c8c9",x"c904",x"c93f",x"c97a",x"c9b5",x"c9f0",x"ca2b",x"ca65",x"ca9f",x"cad9",x"cb13",x"cb4d",x"cb86",x"cbbf",x"cbf8",x"cc31",x"cc6a",x"cca3",x"ccdb",x"cd13",x"cd4b",x"cd83",x"cdbb",x"cdf2",x"ce29",x"ce60",x"ce97",x"cece",x"cf05",x"cf3b",x"cf71",x"cfa7",x"cfdd",x"d013",x"d048",x"d07d",x"d0b3",x"d0e7",x"d11c",x"d151",x"d185",x"d1b9",x"d1ed",x"d221",x"d255",x"d288",x"d2bc",x"d2ef",x"d322",x"d355",x"d387",x"d3ba",x"d3ec",x"d41e",x"d450",x"d482",x"d4b3",x"d4e5",x"d516",x"d547",x"d578",x"d5a8",x"d5d9",x"d609",x"d639",x"d669",x"d699",x"d6c9",x"d6f8",x"d728",x"d757",x"d786",x"d7b4",x"d7e3",x"d811",x"d840",x"d86e",x"d89c",x"d8c9",x"d8f7",x"d924",x"d952",x"d97f",x"d9ac",x"d9d8",x"da05",x"da31",x"da5d",x"da89",x"dab5",x"dae1",x"db0d",x"db38",x"db63",x"db8e",x"dbb9",x"dbe4",x"dc0f",x"dc39",x"dc63",x"dc8d",x"dcb7",x"dce1",x"dd0a",x"dd34",x"dd5d",x"dd86",x"ddaf",x"ddd8",x"de01",x"de29",x"de51",x"de79",x"dea1",x"dec9",x"def1",x"df18",x"df40",x"df67",x"df8e",x"dfb5",x"dfdc",x"e002",x"e029",x"e04f",x"e075",x"e09b",x"e0c1",x"e0e6",x"e10c",x"e131",x"e156",x"e17b",x"e1a0",x"e1c5",x"e1ea",x"e20e",x"e232",x"e256",x"e27a",x"e29e",x"e2c2",x"e2e5",x"e309",x"e32c",x"e34f",x"e372",x"e395",x"e3b8",x"e3da",x"e3fd",x"e41f",x"e441",x"e463",x"e485",x"e4a6",x"e4c8",x"e4e9",x"e50a",x"e52b",x"e54c",x"e56d",x"e58e",x"e5ae",x"e5cf",x"e5ef",x"e60f",x"e62f",x"e64f",x"e66f",x"e68e",x"e6ae",x"e6cd",x"e6ec",x"e70b",x"e72a",x"e749",x"e768",x"e786",x"e7a4",x"e7c3",x"e7e1",x"e7ff",x"e81d",x"e83a",x"e858",x"e875",x"e893",x"e8b0",x"e8cd",x"e8ea",x"e907",x"e923",x"e940",x"e95c",x"e979",x"e995",x"e9b1",x"e9cd",x"e9e9",x"ea04",x"ea20",x"ea3b",x"ea57",x"ea72",x"ea8d",x"eaa8",x"eac3",x"eade",x"eaf8",x"eb13",x"eb2d",x"eb47",x"eb61",x"eb7b",x"eb95",x"ebaf",x"ebc9",x"ebe2",x"ebfc",x"ec15",x"ec2e",x"ec47",x"ec60",x"ec79",x"ec92",x"ecaa",x"ecc3",x"ecdb",x"ecf4",x"ed0c",x"ed24",x"ed3c",x"ed54",x"ed6b",x"ed83",x"ed9b",x"edb2",x"edc9",x"ede1",x"edf8",x"ee0f",x"ee26",x"ee3c",x"ee53",x"ee6a",x"ee80",x"ee96",x"eead",x"eec3",x"eed9",x"eeef",x"ef05",x"ef1a",x"ef30",x"ef46",x"ef5b",x"ef70",x"ef86",x"ef9b",x"efb0",x"efc5",x"efda",x"efee",x"f003",x"f018",x"f02c",x"f040",x"f055",x"f069",x"f07d",x"f091",x"f0a5",x"f0b9",x"f0cc",x"f0e0",x"f0f3",x"f107",x"f11a",x"f12e",x"f141",x"f154",x"f167",x"f17a",x"f18c",x"f19f",x"f1b2",x"f1c4",x"f1d7",x"f1e9",x"f1fb",x"f20d",x"f220",x"f232",x"f243",x"f255",x"f267",x"f279",x"f28a",x"f29c",x"f2ad",x"f2be",x"f2d0",x"f2e1",x"f2f2",x"f303",x"f314",x"f325",x"f335",x"f346",x"f357",x"f367",x"f378",x"f388",x"f398",x"f3a8",x"f3b8",x"f3c9",x"f3d8",x"f3e8",x"f3f8",x"f408",x"f418",x"f427",x"f437",x"f446",x"f455",x"f465",x"f474",x"f483",x"f492",x"f4a1",x"f4b0",x"f4bf",x"f4cd",x"f4dc",x"f4eb",x"f4f9",x"f508",x"f516",x"f525",x"f533",x"f541",x"f54f",x"f55d",x"f56b",x"f579",x"f587",x"f595",x"f5a2",x"f5b0",x"f5be",x"f5cb",x"f5d8",x"f5e6",x"f5f3",x"f600",x"f60e",x"f61b",x"f628",x"f635",x"f642",x"f64e",x"f65b",x"f668",x"f675",x"f681",x"f68e",x"f69a",x"f6a7",x"f6b3",x"f6bf",x"f6cc",x"f6d8",x"f6e4",x"f6f0",x"f6fc",x"f708",x"f714",x"f71f",x"f72b",x"f737",x"f743",x"f74e",x"f75a",x"f765",x"f771",x"f77c",x"f787",x"f792",x"f79e",x"f7a9",x"f7b4",x"f7bf",x"f7ca",x"f7d5",x"f7df",x"f7ea",x"f7f5",x"f800",x"f80a",x"f815",x"f81f",x"f82a",x"f834",x"f83f",x"f849",x"f853",x"f85d",x"f868",x"f872",x"f87c",x"f886",x"f890",x"f89a",x"f8a3",x"f8ad",x"f8b7",x"f8c1",x"f8ca",x"f8d4",x"f8de",x"f8e7",x"f8f1",x"f8fa",x"f903",x"f90d",x"f916",x"f91f",x"f928",x"f931",x"f93b",x"f944",x"f94d",x"f955",x"f95e",x"f967",x"f970",x"f979",x"f982",x"f98a",x"f993",x"f99b",x"f9a4",x"f9ac",x"f9b5",x"f9bd",x"f9c6",x"f9ce",x"f9d6",x"f9df",x"f9e7",x"f9ef",x"f9f7",x"f9ff",x"fa07",x"fa0f",x"fa17",x"fa1f",x"fa27",x"fa2f",x"fa37",x"fa3e",x"fa46",x"fa4e",x"fa55",x"fa5d",x"fa65",x"fa6c",x"fa74",x"fa7b",x"fa82",x"fa8a",x"fa91",x"fa98",x"faa0",x"faa7",x"faae",x"fab5",x"fabc",x"fac3",x"faca",x"fad1",x"fad8",x"fadf",x"fae6",x"faed",x"faf4",x"fafb",x"fb01",x"fb08",x"fb0f",x"fb15",x"fb1c",x"fb23",x"fb29",x"fb30",x"fb36",x"fb3d",x"fb43",x"fb49",x"fb50",x"fb56",x"fb5c",x"fb62",x"fb69",x"fb6f",x"fb75",x"fb7b",x"fb81",x"fb87",x"fb8d",x"fb93",x"fb99",x"fb9f",x"fba5",x"fbab",x"fbb1",x"fbb7",x"fbbc",x"fbc2",x"fbc8",x"fbce",x"fbd3",x"fbd9",x"fbde",x"fbe4",x"fbea",x"fbef",x"fbf5",x"fbfa",x"fbff",x"fc05",x"fc0a",x"fc10",x"fc15",x"fc1a",x"fc1f",x"fc25",x"fc2a",x"fc2f",x"fc34",x"fc39",x"fc3e",x"fc43",x"fc49",x"fc4e",x"fc53",x"fc58",x"fc5c",x"fc61",x"fc66",x"fc6b",x"fc70",x"fc75",x"fc7a",x"fc7e",x"fc83",x"fc88",x"fc8c",x"fc91",x"fc96",x"fc9a",x"fc9f",x"fca4",x"fca8",x"fcad",x"fcb1",x"fcb6",x"fcba",x"fcbf",x"fcc3",x"fcc7",x"fccc",x"fcd0",x"fcd4",x"fcd9",x"fcdd",x"fce1",x"fce5",x"fcea",x"fcee",x"fcf2",x"fcf6",x"fcfa",x"fcfe",x"fd02",x"fd06",x"fd0a",x"fd0e",x"fd12",x"fd16",x"fd1a",x"fd1e",x"fd22",x"fd26",x"fd2a",x"fd2e",x"fd32",x"fd35",x"fd39",x"fd3d",x"fd41",x"fd44",x"fd48",x"fd4c",x"fd4f",x"fd53",x"fd57",x"fd5a",x"fd5e",x"fd61",x"fd65",x"fd69",x"fd6c",x"fd70",x"fd73",x"fd77",x"fd7a",x"fd7d",x"fd81",x"fd84",x"fd88",x"fd8b",x"fd8e",x"fd92",x"fd95",x"fd98",x"fd9b",x"fd9f",x"fda2",x"fda5",x"fda8",x"fdab",x"fdaf",x"fdb2",x"fdb5",x"fdb8",x"fdbb",x"fdbe",x"fdc1",x"fdc4",x"fdc7",x"fdca",x"fdcd",x"fdd0",x"fdd3",x"fdd6",x"fdd9",x"fddc",x"fddf",x"fde2",x"fde5",x"fde8",x"fdeb",x"fded",x"fdf0",x"fdf3",x"fdf6",x"fdf9",x"fdfb",x"fdfe",x"fe01",x"fe03",x"fe06",x"fe09",x"fe0c",x"fe0e",x"fe11",x"fe13",x"fe16",x"fe19",x"fe1b",x"fe1e",x"fe20",x"fe23",x"fe25",x"fe28",x"fe2b",x"fe2d",x"fe2f",x"fe32",x"fe34",x"fe37",x"fe39",x"fe3c",x"fe3e",x"fe40",x"fe43",x"fe45",x"fe48",x"fe4a",x"fe4c",x"fe4f",x"fe51",x"fe53",x"fe55",x"fe58",x"fe5a",x"fe5c",x"fe5e",x"fe61",x"fe63",x"fe65",x"fe67",x"fe69",x"fe6c",x"fe6e",x"fe70",x"fe72",x"fe74",x"fe76",x"fe78",x"fe7a",x"fe7c",x"fe7f",x"fe81",x"fe83",x"fe85",x"fe87",x"fe89",x"fe8b",x"fe8d",x"fe8f",x"fe91",x"fe93",x"fe95",x"fe96",x"fe98",x"fe9a",x"fe9c",x"fe9e",x"fea0",x"fea2",x"fea4",x"fea6",x"fea7",x"fea9",x"feab",x"fead",x"feaf",x"feb0",x"feb2",x"feb4",x"feb6",x"feb8",x"feb9",x"febb",x"febd",x"febe",x"fec0",x"fec2",x"fec4",x"fec5",x"fec7",x"fec9",x"feca",x"fecc",x"fece",x"fecf",x"fed1",x"fed2",x"fed4",x"fed6",x"fed7",x"fed9",x"feda",x"fedc",x"fedd",x"fedf",x"fee1",x"fee2",x"fee4",x"fee5",x"fee7",x"fee8",x"feea",x"feeb",x"feed",x"feee",x"fef0",x"fef1",x"fef2",x"fef4",x"fef5",x"fef7",x"fef8",x"fefa",x"fefb",x"fefc",x"fefe",x"feff",x"ff00",x"ff02",x"ff03",x"ff04",x"ff06",x"ff07",x"ff08",x"ff0a",x"ff0b",x"ff0c",x"ff0e",x"ff0f",x"ff10",x"ff12",x"ff13",x"ff14",x"ff15",x"ff17",x"ff18",x"ff19",x"ff1a",x"ff1c",x"ff1d",x"ff1e",x"ff1f",x"ff20",x"ff22",x"ff23",x"ff24",x"ff25",x"ff26",x"ff27",x"ff29",x"ff2a",x"ff2b",x"ff2c",x"ff2d",x"ff2e",x"ff2f",x"ff30",x"ff32",x"ff33",x"ff34",x"ff35",x"ff36",x"ff37",x"ff38",x"ff39",x"ff3a",x"ff3b",x"ff3c",x"ff3d",x"ff3e",x"ff3f",x"ff40",x"ff41",x"ff42",x"ff44",x"ff45",x"ff46",x"ff47",x"ff47",x"ff48",x"ff49",x"ff4a",x"ff4b",x"ff4c",x"ff4d",x"ff4e",x"ff4f",x"ff50",x"ff51",x"ff52",x"ff53",x"ff54",x"ff55",x"ff56",x"ff57",x"ff58",x"ff58",x"ff59",x"ff5a",x"ff5b",x"ff5c",x"ff5d",x"ff5e",x"ff5f",x"ff5f",x"ff60",x"ff61",x"ff62",x"ff63",x"ff64",x"ff64",x"ff65",x"ff66",x"ff67",x"ff68",x"ff69",x"ff69",x"ff6a",x"ff6b",x"ff6c",x"ff6d",x"ff6d",x"ff6e",x"ff6f",x"ff70",x"ff70",x"ff71",x"ff72",x"ff73",x"ff73",x"ff74",x"ff75",x"ff76",x"ff76",x"ff77",x"ff78",x"ff79",x"ff79",x"ff7a",x"ff7b",x"ff7c",x"ff7c",x"ff7d",x"ff7e",x"ff7e",x"ff7f",x"ff80",x"ff80",x"ff81",x"ff82",x"ff82",x"ff83",x"ff84",x"ff84",x"ff85",x"ff86",x"ff86",x"ff87",x"ff88",x"ff88",x"ff89",x"ff8a",x"ff8a",x"ff8b",x"ff8b",x"ff8c",x"ff8d",x"ff8d",x"ff8e",x"ff8f",x"ff8f",x"ff90",x"ff90",x"ff91",x"ff91",x"ff92",x"ff93",x"ff93",x"ff94",x"ff94",x"ff95",x"ff96",x"ff96",x"ff97",x"ff97",x"ff98",x"ff98",x"ff99",x"ff99",x"ff9a",x"ff9b",x"ff9b",x"ff9c",x"ff9c",x"ff9d",x"ff9d",x"ff9e",x"ff9e",x"ff9f",x"ff9f",x"ffa0",x"ffa0",x"ffa1",x"ffa1",x"ffa2",x"ffa2",x"ffa3",x"ffa3",x"ffa4",x"ffa4",x"ffa5",x"ffa5",x"ffa6",x"ffa6",x"ffa7",x"ffa7",x"ffa8",x"ffa8",x"ffa9",x"ffa9",x"ffaa",x"ffaa",x"ffaa",x"ffab",x"ffab",x"ffac",x"ffac",x"ffad",x"ffad",x"ffae",x"ffae",x"ffae",x"ffaf",x"ffaf",x"ffb0",x"ffb0",x"ffb1",x"ffb1",x"ffb1",x"ffb2",x"ffb2",x"ffb3",x"ffb3",x"ffb4",x"ffb4",x"ffb4",x"ffb5",x"ffb5",x"ffb6",x"ffb6",x"ffb6",x"ffb7",x"ffb7",x"ffb7",x"ffb8",x"ffb8",x"ffb9",x"ffb9",x"ffb9",x"ffba",x"ffba",x"ffbb",x"ffbb",x"ffbb",x"ffbc",x"ffbc",x"ffbc",x"ffbd",x"ffbd",x"ffbd",x"ffbe",x"ffbe",x"ffbe",x"ffbf",x"ffbf",x"ffc0",x"ffc0",x"ffc0",x"ffc1",x"ffc1",x"ffc1",x"ffc2",x"ffc2",x"ffc2",x"ffc3",x"ffc3",x"ffc3",x"ffc4",x"ffc4",x"ffc4",x"ffc4",x"ffc5",x"ffc5",x"ffc5",x"ffc6",x"ffc6",x"ffc6",x"ffc7",x"ffc7",x"ffc7",x"ffc8",x"ffc8",x"ffc8",x"ffc8",x"ffc9",x"ffc9",x"ffc9",x"ffca",x"ffca",x"ffca",x"ffca",x"ffcb",x"ffcb",x"ffcb",x"ffcc",x"ffcc",x"ffcc",x"ffcc",x"ffcd",x"ffcd",x"ffcd",x"ffce",x"ffce",x"ffce",x"ffce",x"ffcf",x"ffcf",x"ffcf",x"ffcf",x"ffd0",x"ffd0",x"ffd0",x"ffd0",x"ffd1",x"ffd1",x"ffd1",x"ffd1",x"ffd2",x"ffd2",x"ffd2",x"ffd2",x"ffd3",x"ffd3",x"ffd3",x"ffd3",x"ffd4",x"ffd4",x"ffd4",x"ffd4",x"ffd4",x"ffd5",x"ffd5",x"ffd5",x"ffd5",x"ffd6",x"ffd6",x"ffd6",x"ffd6",x"ffd7",x"ffd7",x"ffd7",x"ffd7",x"ffd7",x"ffd8",x"ffd8",x"ffd8",x"ffd8",x"ffd8",x"ffd9",x"ffd9",x"ffd9",x"ffd9",x"ffd9",x"ffda",x"ffda",x"ffda",x"ffda",x"ffda",x"ffdb",x"ffdb",x"ffdb",x"ffdb",x"ffdb",x"ffdc",x"ffdc",x"ffdc",x"ffdc",x"ffdc",x"ffdd",x"ffdd",x"ffdd",x"ffdd",x"ffdd",x"ffde",x"ffde",x"ffde",x"ffde",x"ffde",x"ffde",x"ffdf",x"ffdf",x"ffdf",x"ffdf",x"ffdf",x"ffdf",x"ffe0",x"ffe0",x"ffe0",x"ffe0",x"ffe0",x"ffe0",x"ffe1",x"ffe1",x"ffe1",x"ffe1",x"ffe1",x"ffe1",x"ffe2",x"ffe2",x"ffe2",x"ffe2",x"ffe2",x"ffe2",x"ffe3",x"ffe3",x"ffe3",x"ffe3",x"ffe3",x"ffe3",x"ffe4",x"ffe4",x"ffe4",x"ffe4",x"ffe4",x"ffe4",x"ffe4",x"ffe5",x"ffe5",x"ffe5",x"ffe5",x"ffe5",x"ffe5",x"ffe5",x"ffe6",x"ffe6",x"ffe6",x"ffe6",x"ffe6",x"ffe6",x"ffe6",x"ffe6",x"ffe7",x"ffe7",x"ffe7",x"ffe7",x"ffe7",x"ffe7",x"ffe7",x"ffe8",x"ffe8",x"ffe8",x"ffe8",x"ffe8",x"ffe8",x"ffe8",x"ffe8",x"ffe9",x"ffe9",x"ffe9",x"ffe9",x"ffe9",x"ffe9",x"ffe9",x"ffe9",x"ffea",x"ffea",x"ffea",x"ffea",x"ffea",x"ffea",x"ffea",x"ffea",x"ffea",x"ffeb",x"ffeb",x"ffeb",x"ffeb",x"ffeb",x"ffeb",x"ffeb",x"ffeb",x"ffeb",x"ffec",x"ffec",x"ffec",x"ffec",x"ffec",x"ffec",x"ffec",x"ffec",x"ffec",x"ffec",x"ffed",x"ffed",x"ffed",x"ffed",x"ffed",x"ffed",x"ffed",x"ffed",x"ffed",x"ffed",x"ffee",x"ffee",x"ffee",x"ffee",x"ffee",x"ffee",x"ffee",x"ffee",x"ffee",x"ffee",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"ffef",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff0",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff1",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff2",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff3",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff4",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff5",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff6",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff7",x"fff8",x"fff8",x"fff8",x"fff9",x"fff9",x"fff9",x"fffa",x"fffa",x"fffa",x"fffa",x"fffa",x"fffb",x"fffb",x"fffb",x"fffb",x"fffb",x"fffc",x"fffc",x"fffc",x"fffc",x"fffc",x"fffc",x"fffd",x"fffd",x"fffd",x"fffe",x"fffe",x"fffe",x"fffe");
    signal ind, dec, decimal_32, ent_32 : integer := 0;
begin
    
    process (clk) begin
        if rising_edge(clk) then
            decimal_32 <=  conv_integer(x"0000" & Y(15 downto 0));
            ent_32 <= conv_integer(Y(31 downto 16));
        end if;    
    end process;
    
    process (clk) begin
        if rising_edge(clk) then
            if ( Y(31 downto 16) < -10 ) then 
                dec <= decimal_32/9855;
            elsif ( Y(31 downto 16) < -9 ) then 
                dec <= decimal_32/2815;
            elsif ( Y(31 downto 16) < 9 ) then 
                dec <= decimal_32/351;
            elsif ( Y(31 downto 16) < 10 ) then 
                dec <= decimal_32/2815;
            else 
                dec <= decimal_32/9855;
            end if;
        end if;
    end process;
    
    process (clk) begin
        if rising_edge(clk) then
            if ( Y(31 downto 16) < -10 ) then 
                ind <= dec;
            elsif ( Y(31 downto 16) < -9 ) then 
                ind <= 7 + dec;
            elsif ( Y(31 downto 16) < 9 ) then 
                ind <= 1704+(ent_32*186)+dec;
            elsif ( Y(31 downto 16) < 10 ) then 
                ind <= 1705+(ent_32*186)+dec;
            else
                ind <= 1728+(ent_32*186)+dec; 
            end if;
        end if;
    end process;
    
    process (clk) begin
        if rising_edge(clk) then
            if (Y(31 downto 16) < -11) then O <= x"00000000";
            elsif (Y(31 downto 16) > 11) then O <= x"0000FFFF";
            else
             O <= x"0000" & sigmoid_val(ind);
            end if; 
        end if;
    end process;
         
end Behavioral;
